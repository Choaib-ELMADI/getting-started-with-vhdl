entity wait_on_wait_until_tb is
end entity;

architecture sim of wait_on_wait_until_tb is
begin

    process is
    begin

        
        

    end process;

end architecture;
