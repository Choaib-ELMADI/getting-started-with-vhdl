entity wait_tb is
end entity;

architecture sim of wait_tb is
begin:

    wait;   -- Indefinitely stop the program execution

end architecture;
