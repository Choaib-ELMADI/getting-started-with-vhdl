entity report_tb is
end entity;

architecture sim of report_tb is
begin:

    report "Hello, World!"; -- Print messages on the simulator console
    wait;

end architecture;
