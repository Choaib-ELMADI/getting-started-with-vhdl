entity tb_0_hello_world is
end entity;

architecture sim of tb_0_hello_world is
begin

    process is
    begin

        report "Hello, World! YEAAAH";
        wait;

    end process;

end architecture;
